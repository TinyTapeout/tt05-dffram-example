VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM32
  CLASS BLOCK ;
  FOREIGN RAM32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 401.580 BY 136.000 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 17.720 401.580 18.320 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 29.960 401.580 30.560 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 42.200 401.580 42.800 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 54.440 401.580 55.040 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 66.680 401.580 67.280 ;
    END
  END A0[4]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 399.580 78.920 401.580 79.520 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 7.910 134.000 8.190 136.000 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 134.000 132.390 136.000 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 144.530 134.000 144.810 136.000 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 156.950 134.000 157.230 136.000 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 169.370 134.000 169.650 136.000 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 181.790 134.000 182.070 136.000 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 194.210 134.000 194.490 136.000 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 206.630 134.000 206.910 136.000 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 134.000 219.330 136.000 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 231.470 134.000 231.750 136.000 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 243.890 134.000 244.170 136.000 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 20.330 134.000 20.610 136.000 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 256.310 134.000 256.590 136.000 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 268.730 134.000 269.010 136.000 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 281.150 134.000 281.430 136.000 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 293.570 134.000 293.850 136.000 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 305.990 134.000 306.270 136.000 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 318.410 134.000 318.690 136.000 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 330.830 134.000 331.110 136.000 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 343.250 134.000 343.530 136.000 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 355.670 134.000 355.950 136.000 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 368.090 134.000 368.370 136.000 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 32.750 134.000 33.030 136.000 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 380.510 134.000 380.790 136.000 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 134.000 393.210 136.000 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 134.000 45.450 136.000 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 57.590 134.000 57.870 136.000 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 70.010 134.000 70.290 136.000 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 82.430 134.000 82.710 136.000 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 94.850 134.000 95.130 136.000 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 107.270 134.000 107.550 136.000 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 119.690 134.000 119.970 136.000 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 5.480 401.580 6.080 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.580 2.480 23.180 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.180 2.480 176.780 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.780 2.480 330.380 133.520 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.520 21.870 399.060 23.470 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 133.520 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.520 18.570 399.060 20.170 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 91.160 401.580 91.760 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 103.400 401.580 104.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 115.640 401.580 116.240 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 127.880 401.580 128.480 ;
    END
  END WE0[3]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 398.820 133.365 ;
      LAYER met1 ;
        RECT 2.760 0.040 398.820 135.960 ;
      LAYER met2 ;
        RECT 3.310 133.720 7.630 135.990 ;
        RECT 8.470 133.720 20.050 135.990 ;
        RECT 20.890 133.720 32.470 135.990 ;
        RECT 33.310 133.720 44.890 135.990 ;
        RECT 45.730 133.720 57.310 135.990 ;
        RECT 58.150 133.720 69.730 135.990 ;
        RECT 70.570 133.720 82.150 135.990 ;
        RECT 82.990 133.720 94.570 135.990 ;
        RECT 95.410 133.720 106.990 135.990 ;
        RECT 107.830 133.720 119.410 135.990 ;
        RECT 120.250 133.720 131.830 135.990 ;
        RECT 132.670 133.720 144.250 135.990 ;
        RECT 145.090 133.720 156.670 135.990 ;
        RECT 157.510 133.720 169.090 135.990 ;
        RECT 169.930 133.720 181.510 135.990 ;
        RECT 182.350 133.720 193.930 135.990 ;
        RECT 194.770 133.720 206.350 135.990 ;
        RECT 207.190 133.720 218.770 135.990 ;
        RECT 219.610 133.720 231.190 135.990 ;
        RECT 232.030 133.720 243.610 135.990 ;
        RECT 244.450 133.720 256.030 135.990 ;
        RECT 256.870 133.720 268.450 135.990 ;
        RECT 269.290 133.720 280.870 135.990 ;
        RECT 281.710 133.720 293.290 135.990 ;
        RECT 294.130 133.720 305.710 135.990 ;
        RECT 306.550 133.720 318.130 135.990 ;
        RECT 318.970 133.720 330.550 135.990 ;
        RECT 331.390 133.720 342.970 135.990 ;
        RECT 343.810 133.720 355.390 135.990 ;
        RECT 356.230 133.720 367.810 135.990 ;
        RECT 368.650 133.720 380.230 135.990 ;
        RECT 381.070 133.720 392.650 135.990 ;
        RECT 393.490 133.720 397.340 135.990 ;
        RECT 3.310 2.280 397.340 133.720 ;
        RECT 3.310 0.010 7.630 2.280 ;
        RECT 8.470 0.010 20.050 2.280 ;
        RECT 20.890 0.010 32.470 2.280 ;
        RECT 33.310 0.010 44.890 2.280 ;
        RECT 45.730 0.010 57.310 2.280 ;
        RECT 58.150 0.010 69.730 2.280 ;
        RECT 70.570 0.010 82.150 2.280 ;
        RECT 82.990 0.010 94.570 2.280 ;
        RECT 95.410 0.010 106.990 2.280 ;
        RECT 107.830 0.010 119.410 2.280 ;
        RECT 120.250 0.010 131.830 2.280 ;
        RECT 132.670 0.010 144.250 2.280 ;
        RECT 145.090 0.010 156.670 2.280 ;
        RECT 157.510 0.010 169.090 2.280 ;
        RECT 169.930 0.010 181.510 2.280 ;
        RECT 182.350 0.010 193.930 2.280 ;
        RECT 194.770 0.010 206.350 2.280 ;
        RECT 207.190 0.010 218.770 2.280 ;
        RECT 219.610 0.010 231.190 2.280 ;
        RECT 232.030 0.010 243.610 2.280 ;
        RECT 244.450 0.010 256.030 2.280 ;
        RECT 256.870 0.010 268.450 2.280 ;
        RECT 269.290 0.010 280.870 2.280 ;
        RECT 281.710 0.010 293.290 2.280 ;
        RECT 294.130 0.010 305.710 2.280 ;
        RECT 306.550 0.010 318.130 2.280 ;
        RECT 318.970 0.010 330.550 2.280 ;
        RECT 331.390 0.010 342.970 2.280 ;
        RECT 343.810 0.010 355.390 2.280 ;
        RECT 356.230 0.010 367.810 2.280 ;
        RECT 368.650 0.010 380.230 2.280 ;
        RECT 381.070 0.010 392.650 2.280 ;
        RECT 393.490 0.010 397.340 2.280 ;
      LAYER met3 ;
        RECT 3.285 128.880 399.580 135.825 ;
        RECT 3.285 127.480 399.180 128.880 ;
        RECT 3.285 116.640 399.580 127.480 ;
        RECT 3.285 115.240 399.180 116.640 ;
        RECT 3.285 104.400 399.580 115.240 ;
        RECT 3.285 103.000 399.180 104.400 ;
        RECT 3.285 92.160 399.580 103.000 ;
        RECT 3.285 90.760 399.180 92.160 ;
        RECT 3.285 79.920 399.580 90.760 ;
        RECT 3.285 78.520 399.180 79.920 ;
        RECT 3.285 67.680 399.580 78.520 ;
        RECT 3.285 66.280 399.180 67.680 ;
        RECT 3.285 55.440 399.580 66.280 ;
        RECT 3.285 54.040 399.180 55.440 ;
        RECT 3.285 43.200 399.580 54.040 ;
        RECT 3.285 41.800 399.180 43.200 ;
        RECT 3.285 30.960 399.580 41.800 ;
        RECT 3.285 29.560 399.180 30.960 ;
        RECT 3.285 18.720 399.580 29.560 ;
        RECT 3.285 17.320 399.180 18.720 ;
        RECT 3.285 6.480 399.580 17.320 ;
        RECT 3.285 5.080 399.180 6.480 ;
        RECT 3.285 0.175 399.580 5.080 ;
      LAYER met4 ;
        RECT 90.455 6.295 171.480 79.385 ;
        RECT 173.880 6.295 174.780 79.385 ;
        RECT 177.180 6.295 325.080 79.385 ;
        RECT 327.480 6.295 328.380 79.385 ;
        RECT 330.780 6.295 391.625 79.385 ;
  END
END RAM32
END LIBRARY

